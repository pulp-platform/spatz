../src/generated/testharness.sv